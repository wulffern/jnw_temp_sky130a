*TB_SUN_TR_SKY130NM/TB_NCM



*----------------------------------------------------------------
* Include
*----------------------------------------------------------------

.include ../../../../cpdk/ngspice/ideal_circuits.spi


#ifdef Lay
.include ../../../work/lpe/JNW_TEMP_lpe.spi
#else
.include ../../../work/xsch/JNW_TEMP.spice
#endif



*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15
*reltol=1e-4 method=gear

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

.param PERIOD_CLK = 1/50e6

.param PW_CLK = PERIOD_CLK/2

.param TSTART = 10n

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD_1V8  0 pwl 0 0 {TSTART/2} {AVDD}
*VCLK clk 0 dc 0
*VRESET reset 0 dc 0
VCLK clk 0 dc 0 pulse (0 {AVDD} {TSTART} {TRF} {TRF} {PW_CLK} {PERIOD_CLK})
VRESET reset 0 dc {AVDD} pwl {TSTART} {AVDD} {PW_CLK} {AVDD} {PW_CLK*2} 0



*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi
.include ../svinst.spi

*- Fakearoony to get the digital sha included. Never actually included
*#include ../../../rtl/dig.v



.save V(PWM_1V8)
.save v(din)
.save v(xdut.xibps.vr1)
.save v(xdut.xibps.vd1)
.save v(xdut.xibps.vd2)
.save v(xdut.xibp.vd2)
.save v(xdut.xibp.vd1)
.save v(xdut.xibp.vr1)
.save v(xdut.ibps_1u<2>)
.save v(xdut.ibps_1u<1>)
.save v(xdut.ibp_1u<0>)
.save v(xdut.ibp_1u<2>)
.save v(xdut.ibp_1u<3>)
.save v(xdut.ibp_1u<1>) v(CMPO_1V8) v(xdut.vip)
*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
#ifdef Nosweep
.save all
#endif


*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

*- Override the default digital output bridge.
pre_set auto_bridge_d_out =
     + ( ".model auto_dac dac_bridge(out_low = 0.0 out_high = 1.8)"
     +   "auto_bridge%d [ %s ] [ %s ] auto_dac" )


optran 0 0 0 1n 1u 0


set fend = .raw
#ifdef Nosweep
*.option temp=42.5
*.option temp=-40
tran 1n 6u
write {cicname}.raw
#else
foreach vtemp {temperatures}
  option temp=$vtemp
  tran 1n 10u 4u
  write {cicname}_$vtemp$fend
end

#endif

quit


.endc

.end
